.title KiCad schematic
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/LP38693_ADJ_TRANS.lib"
.include "models/PCF1C101MCL1GS_v100.lib"
.include "models/PCF1E100MCL1GS_v100.lib"
XU3 VCC /ADJ /EN /OUT 0 LP38693_ADJ_TRANS
R1 VCC /EN {Ren}
R2 /OUT /ADJ {Radj}
R3 /ADJ 0 {Rref}
XU1 VCC 0 PCF1E100MCL1GS
XU4 /OUT 0 PCF1C101MCL1GS
XU2 VCC 0 C2012X7R2A104K125AA_p
V1 VCC 0 {VIN}
I1 0 /OUT {ILOAD}
XU5 /OUT 0 C2012X7R2A104K125AA_p
.end
